// This logic just worked, I haven't simplified the truth table
module top_module (
    input a,
    input b,
    input c,
    input d,
    output q );//

    assign q = c | b ; // Fix me

endmodule
